module Mux8 (
    input wire [7:0] inputA,
    input wire [7:0] inputB,
    input wire control,

    output reg [7:0] muxed
);
    
endmodule